-- @author EliasDH Team
-- @see https://eliasdh.com
-- @since 01/01/2025